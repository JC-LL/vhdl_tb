-- blah
-- entity
library ieee;
use ieee.std_logic_1164.all;

entity test1 is
   
end;

architecture rtl of test1 is
begin
end rtl;
